5202|0676529|NMB|Barker, Nick
20095|9974948|MPB|Barrow, Mark
20192|1371522|NB|Barry, Nicolas
13816|1172494|LB|Bayley, Lynne
252|0380634|CAB|Blindauer, Claudia
236|9775013|SAFB|Bon, Stefan
7688|0971041|JB|Brannon, Julie
15899|0270199|SB|Brown, Steven
235|9970029|TDHB|Bugg, Tim
232|0070559|GLC|Challis, Gregory L
11297|1074204|ABC|Chaplin, Adrian
12692|1070634|NC|Chmel, Nikola
253|9370232|AJC|Clark, Andrew
264|9871900|GJC|Clarkson, Guy J
11634|0670255|SC|Coles, Stuart
9217|0380711|CC|Corre, Christophe
3470|0674312|GC|Costantini, Giovanni
14929|0070384|JAC|Covington, James
20241|0974163|CDGC|Cunningham, Charlie
18435|1274901|GLD|Davies, Gemma-Louise
9354|038057|GDC|De Calvo, Gillian
250|9573369|RJD|Deeth, Rob
234|0482387|AMD|Dixon, Ann
237|0483339|APD|Dove, Andrew
1419|0670020|DJF|Fox, David
11697|1171759|JG|Geden, Jo
9437|0970074|MIG|Gibson, Matt
13765|1172916|SH|Habershon, Scott
12114|0673019|AH|Habtemariam, Abraha
222|9370782|DMH|Haddleton, David
5780|0770905|RH|Hatton, Ross
3089|0671811|TSJ|Jones, Tim
10974|1071602|JRL|Lewandowski, Jozef
231|0770308|IM|Mackirdy, Ian
244|9671494|JVM|Macpherson, Julie
230|9576089|AM|Marsh, Andrew
9219|0874020|RN|Notman, Rebecca
6860|0871340|PBO|O'Connor, Peter
5806|0871352|RKO|O'Reilly Rachel
14122|1270619|GP|Pattison, Graham
17119|1274179|SP|Perrier, Sebastian
11299|0770882|IP|Prokes, Ivan
233|9471544|AR|Rodger, Alison
249|9876059|PMR|Rodger, Mark
20233|u1374301|DR|Roper, Daniel
243|9470222|JPR|Rourke, Jon
3088|0671901|PJS|Sadler, Peter J
240|9677551|PS|Scott, Peter
241|0370203|MS|Shipman, Mike
11298|0580038|LS|Song, Lijiang
263|0482356|VS|Stavros, Vasilios
260|9170320|PCT|Taylor, Paul
9713|1070530|MT|Tosin, Manuela
225|0483109|AT|Troisi, Alessandro
17621|9678316|SU|Udall, Sharon
256|9172223|PRU|Unwin, Pat
259|0582691|RIW|Walton, Richard
254|0370604|GW|Willey, Gerald
238|9574780|MW|Wills, Martin
20445|0971273|PW|Wilson, Paul
9877234|9877234|JN|Noone, Jason
261|||Everyone
266|||External
9544|8670364|JE|Emmerson, Jane
9407|0970410|EH|Hardiman, Elizabeth
9503|||Hicks, Matthew
12691|||Howarth, Oliver
17618|1071657|CM|Martin, Claire
14971|||Steven Howdle
21396|1473674|PC|Paolo Coppo
21395|1474109|RK|Russ Kitson
